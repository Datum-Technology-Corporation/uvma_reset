// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_RESET_ST_MACROS_SV__
`define __UVME_RESET_ST_MACROS_SV__





`endif // __UVME_RESET_ST_MACROS_SV__
