// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_RESET_ST_TDEFS_SV__
`define __UVMT_RESET_ST_TDEFS_SV__





`endif // __UVMT_RESET_ST_TDEFS_SV__
