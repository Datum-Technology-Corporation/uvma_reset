// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_RESET_ST_CONSTANTS_SV__
`define __UVME_RESET_ST_CONSTANTS_SV__


const int unsigned  uvme_reset_st_rand_pulses_default_num_pulses          =    10;
const int unsigned  uvme_reset_st_rand_pulses_default_min_pulse_duration  =     1;
const int unsigned  uvme_reset_st_rand_pulses_default_max_pulse_duration  =   100;
const int unsigned  uvme_reset_st_rand_pulses_default_min_pulse_gap       =   100;
const int unsigned  uvme_reset_st_rand_pulses_default_max_pulse_gap       = 1_000;


`endif // __UVME_RESET_ST_CONSTANTS_SV__
