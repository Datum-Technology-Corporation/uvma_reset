// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_RESET_IF_CHKR_SV__
`define __UVMA_RESET_IF_CHKR_SV__


/**
 * Encapsulates assertions targeting uvma_reset_if.
 */
module uvma_reset_if_chkr(
   uvma_reset_if  reset_if
);
   
   // TODO Add assertions to uvma_reset_if_chkr
   
endmodule : uvma_reset_if_chkr


`endif // __UVMA_RESET_IF_CHKR_SV__
